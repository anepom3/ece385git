// This file is for the NZP register!
