// This file is for the BEN register!
