// This is the file for the SR1MUX!
