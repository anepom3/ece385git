// We'll create the MDR module here!
