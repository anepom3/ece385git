// This file is for the REGFILE module!
