// This file is for the ALU module.
