// We'll create the MAR module here.
// This is just a 16-bit register.
