module Shooter ();
  
endmodule // Shooter
