// TODO we'l make a datapath module here!
// This will be used to connect all the modules together.
// PC (Program Counter) Package: PC, PCMUX, '+1', GatePC
// MDR Package: MDR, GateMDR
// MAR Package: MAR, GateMAR
// IR Package: IR
// 
