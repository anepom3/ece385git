// This is the file for the SR2MUX!
