module Barrier ( input level_sel,
                 output logic [0:14][0:19] barrier // include [0:1] --> ...[0:19][0:1] barrier
  );

  always_comb begin

    case (level_sel)
      0:
      barrier <=
        '{
        '{1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
        '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}
        };
      1:
        barrier <=
          '{
          '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
          '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
          '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
          '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
          '{0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0},
          '{0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0},
          '{0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0},
          '{0,0,0,1,0,0,0,1,0,0,0,0,0,0,0,0,1,0,0,0},
          '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
          '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
          '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
          '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
          '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
          '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
          '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}
          };
      default:
        barrier <=
          '{
          '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
          '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
          '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
          '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
          '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
          '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
          '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
          '{0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0},
          '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
          '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
          '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
          '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
          '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
          '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
          '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}
          };
    endcase
  end
endmodule // barrier
