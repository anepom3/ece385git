// We'll create the program counter module here!
