// This is the file for the ADDR1MUX!
