module cla_4bit
(
    input   logic[3:0]     A,
    input   logic[3:0]     B,
    output  logic[3:0]     Sum,
    output  logic           CO,
	 output  logic          Pg,
	 output  logic          Gg
);

















endmodule
