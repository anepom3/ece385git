// We'll create the MDR module here!
// This is just a 16-bit register.
