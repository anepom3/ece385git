// This file will be for the GatePC, GateMAR, GateMDR, and GateALU tristate
// buffers. (It will actually just be a 5-to-1 MUX, 5th being 16'hxxxx)
