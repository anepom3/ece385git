// We'll create the IR file here!
// This is just a 16-bit register.
