// TODO we'l make a datapath module here!
