// This is the file for the DRMUX!
