// lab9_soc.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module lab9_soc (
		output wire [31:0] aes_export_export_data,                        //                             aes_export.export_data
		input  wire        clk_clk,                                       //                                    clk.clk
		output wire        nios2_gen2_0_custom_instruction_master_readra, // nios2_gen2_0_custom_instruction_master.readra
		input  wire        reset_reset_n,                                 //                                  reset.reset_n
		output wire        sdram_clk_clk,                                 //                              sdram_clk.clk
		output wire [12:0] sdram_wire_addr,                               //                             sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                                 //                                       .ba
		output wire        sdram_wire_cas_n,                              //                                       .cas_n
		output wire        sdram_wire_cke,                                //                                       .cke
		output wire        sdram_wire_cs_n,                               //                                       .cs_n
		inout  wire [15:0] sdram_wire_dq,                                 //                                       .dq
		output wire [1:0]  sdram_wire_dqm,                                //                                       .dqm
		output wire        sdram_wire_ras_n,                              //                                       .ras_n
		output wire        sdram_wire_we_n                                //                                       .we_n
	);

	wire         sdram_pll_c0_clk;                                             // SDRAM_PLL:c0 -> [SDRAM:clk, mm_interconnect_0:SDRAM_PLL_c0_clk, rst_controller_001:clk]
	wire  [31:0] nios2_data_master_readdata;                                   // mm_interconnect_0:NIOS2_data_master_readdata -> NIOS2:d_readdata
	wire         nios2_data_master_waitrequest;                                // mm_interconnect_0:NIOS2_data_master_waitrequest -> NIOS2:d_waitrequest
	wire         nios2_data_master_debugaccess;                                // NIOS2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOS2_data_master_debugaccess
	wire  [27:0] nios2_data_master_address;                                    // NIOS2:d_address -> mm_interconnect_0:NIOS2_data_master_address
	wire   [3:0] nios2_data_master_byteenable;                                 // NIOS2:d_byteenable -> mm_interconnect_0:NIOS2_data_master_byteenable
	wire         nios2_data_master_read;                                       // NIOS2:d_read -> mm_interconnect_0:NIOS2_data_master_read
	wire         nios2_data_master_write;                                      // NIOS2:d_write -> mm_interconnect_0:NIOS2_data_master_write
	wire  [31:0] nios2_data_master_writedata;                                  // NIOS2:d_writedata -> mm_interconnect_0:NIOS2_data_master_writedata
	wire  [31:0] nios2_instruction_master_readdata;                            // mm_interconnect_0:NIOS2_instruction_master_readdata -> NIOS2:i_readdata
	wire         nios2_instruction_master_waitrequest;                         // mm_interconnect_0:NIOS2_instruction_master_waitrequest -> NIOS2:i_waitrequest
	wire  [27:0] nios2_instruction_master_address;                             // NIOS2:i_address -> mm_interconnect_0:NIOS2_instruction_master_address
	wire         nios2_instruction_master_read;                                // NIOS2:i_read -> mm_interconnect_0:NIOS2_instruction_master_read
	wire         mm_interconnect_0_aes_decryption_core_0_aes_slave_chipselect; // mm_interconnect_0:AES_Decryption_Core_0_AES_Slave_chipselect -> AES_Decryption_Core_0:AVL_CS
	wire  [31:0] mm_interconnect_0_aes_decryption_core_0_aes_slave_readdata;   // AES_Decryption_Core_0:AVL_READDATA -> mm_interconnect_0:AES_Decryption_Core_0_AES_Slave_readdata
	wire   [3:0] mm_interconnect_0_aes_decryption_core_0_aes_slave_address;    // mm_interconnect_0:AES_Decryption_Core_0_AES_Slave_address -> AES_Decryption_Core_0:AVL_ADDR
	wire         mm_interconnect_0_aes_decryption_core_0_aes_slave_read;       // mm_interconnect_0:AES_Decryption_Core_0_AES_Slave_read -> AES_Decryption_Core_0:AVL_READ
	wire   [3:0] mm_interconnect_0_aes_decryption_core_0_aes_slave_byteenable; // mm_interconnect_0:AES_Decryption_Core_0_AES_Slave_byteenable -> AES_Decryption_Core_0:AVL_BYTE_EN
	wire         mm_interconnect_0_aes_decryption_core_0_aes_slave_write;      // mm_interconnect_0:AES_Decryption_Core_0_AES_Slave_write -> AES_Decryption_Core_0:AVL_WRITE
	wire  [31:0] mm_interconnect_0_aes_decryption_core_0_aes_slave_writedata;  // mm_interconnect_0:AES_Decryption_Core_0_AES_Slave_writedata -> AES_Decryption_Core_0:AVL_WRITEDATA
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;     // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_chipselect -> JTAG_UART:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;       // JTAG_UART:av_readdata -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;    // JTAG_UART:av_waitrequest -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;        // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_address -> JTAG_UART:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;           // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_read -> JTAG_UART:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;          // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_write -> JTAG_UART:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;      // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_writedata -> JTAG_UART:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_sysid_control_slave_readdata;         // NIOS2_SYSID:readdata -> mm_interconnect_0:NIOS2_SYSID_control_slave_readdata
	wire   [0:0] mm_interconnect_0_nios2_sysid_control_slave_address;          // mm_interconnect_0:NIOS2_SYSID_control_slave_address -> NIOS2_SYSID:address
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_readdata;             // NIOS2:debug_mem_slave_readdata -> mm_interconnect_0:NIOS2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_debug_mem_slave_waitrequest;          // NIOS2:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOS2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_debug_mem_slave_debugaccess;          // mm_interconnect_0:NIOS2_debug_mem_slave_debugaccess -> NIOS2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_debug_mem_slave_address;              // mm_interconnect_0:NIOS2_debug_mem_slave_address -> NIOS2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_debug_mem_slave_read;                 // mm_interconnect_0:NIOS2_debug_mem_slave_read -> NIOS2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_debug_mem_slave_byteenable;           // mm_interconnect_0:NIOS2_debug_mem_slave_byteenable -> NIOS2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_debug_mem_slave_write;                // mm_interconnect_0:NIOS2_debug_mem_slave_write -> NIOS2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_writedata;            // mm_interconnect_0:NIOS2_debug_mem_slave_writedata -> NIOS2:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_readdata;               // SDRAM_PLL:readdata -> mm_interconnect_0:SDRAM_PLL_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_sdram_pll_pll_slave_address;                // mm_interconnect_0:SDRAM_PLL_pll_slave_address -> SDRAM_PLL:address
	wire         mm_interconnect_0_sdram_pll_pll_slave_read;                   // mm_interconnect_0:SDRAM_PLL_pll_slave_read -> SDRAM_PLL:read
	wire         mm_interconnect_0_sdram_pll_pll_slave_write;                  // mm_interconnect_0:SDRAM_PLL_pll_slave_write -> SDRAM_PLL:write
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_writedata;              // mm_interconnect_0:SDRAM_PLL_pll_slave_writedata -> SDRAM_PLL:writedata
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;                // mm_interconnect_0:ONCHIP_MEMORY_s1_chipselect -> ONCHIP_MEMORY:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;                  // ONCHIP_MEMORY:readdata -> mm_interconnect_0:ONCHIP_MEMORY_s1_readdata
	wire   [1:0] mm_interconnect_0_onchip_memory_s1_address;                   // mm_interconnect_0:ONCHIP_MEMORY_s1_address -> ONCHIP_MEMORY:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;                // mm_interconnect_0:ONCHIP_MEMORY_s1_byteenable -> ONCHIP_MEMORY:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                     // mm_interconnect_0:ONCHIP_MEMORY_s1_write -> ONCHIP_MEMORY:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;                 // mm_interconnect_0:ONCHIP_MEMORY_s1_writedata -> ONCHIP_MEMORY:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                     // mm_interconnect_0:ONCHIP_MEMORY_s1_clken -> ONCHIP_MEMORY:clken
	wire         mm_interconnect_0_sdram_s1_chipselect;                        // mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                          // SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                       // SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                           // mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                              // mm_interconnect_0:SDRAM_s1_read -> SDRAM:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                        // mm_interconnect_0:SDRAM_s1_byteenable -> SDRAM:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                     // SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                             // mm_interconnect_0:SDRAM_s1_write -> SDRAM:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                         // mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	wire         irq_mapper_receiver0_irq;                                     // JTAG_UART:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_irq_irq;                                                // irq_mapper:sender_irq -> NIOS2:irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [AES_Decryption_Core_0:RESET, JTAG_UART:rst_n, NIOS2:reset_n, NIOS2_SYSID:reset_n, ONCHIP_MEMORY:reset, SDRAM_PLL:reset, irq_mapper:reset, mm_interconnect_0:NIOS2_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [NIOS2:reset_req, ONCHIP_MEMORY:reset_req, rst_translator:reset_req_in]
	wire         nios2_debug_reset_request_reset;                              // NIOS2:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                           // rst_controller_001:reset_out -> [SDRAM:reset_n, mm_interconnect_0:SDRAM_reset_reset_bridge_in_reset_reset]

	avalon_aes_interface aes_decryption_core_0 (
		.CLK           (clk_clk),                                                      //         CLK.clk
		.RESET         (rst_controller_reset_out_reset),                               //       RESET.reset
		.AVL_CS        (mm_interconnect_0_aes_decryption_core_0_aes_slave_chipselect), //   AES_Slave.chipselect
		.AVL_BYTE_EN   (mm_interconnect_0_aes_decryption_core_0_aes_slave_byteenable), //            .byteenable
		.AVL_ADDR      (mm_interconnect_0_aes_decryption_core_0_aes_slave_address),    //            .address
		.AVL_WRITEDATA (mm_interconnect_0_aes_decryption_core_0_aes_slave_writedata),  //            .writedata
		.AVL_READDATA  (mm_interconnect_0_aes_decryption_core_0_aes_slave_readdata),   //            .readdata
		.AVL_WRITE     (mm_interconnect_0_aes_decryption_core_0_aes_slave_write),      //            .write
		.AVL_READ      (mm_interconnect_0_aes_decryption_core_0_aes_slave_read),       //            .read
		.EXPORT_DATA   (aes_export_export_data)                                        // EXPORT_DATA.export_data
	);

	lab9_soc_JTAG_UART jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	lab9_soc_NIOS2 nios2 (
		.clk                                 (clk_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (nios2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       (nios2_gen2_0_custom_instruction_master_readra)        // custom_instruction_master.readra
	);

	lab9_soc_NIOS2_SYSID nios2_sysid (
		.clock    (clk_clk),                                              //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                      //         reset.reset_n
		.readdata (mm_interconnect_0_nios2_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_nios2_sysid_control_slave_address)   //              .address
	);

	lab9_soc_ONCHIP_MEMORY onchip_memory (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),            //       .reset_req
		.freeze     (1'b0)                                           // (terminated)
	);

	lab9_soc_SDRAM sdram (
		.clk            (sdram_pll_c0_clk),                         //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	lab9_soc_SDRAM_PLL sdram_pll (
		.clk                (clk_clk),                                         //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset),                  // inclk_interface_reset.reset
		.read               (mm_interconnect_0_sdram_pll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_sdram_pll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_sdram_pll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_sdram_pll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_sdram_pll_pll_slave_writedata), //                      .writedata
		.c0                 (sdram_pll_c0_clk),                                //                    c0.clk
		.c1                 (sdram_clk_clk),                                   //                    c1.clk
		.scandone           (),                                                //           (terminated)
		.scandataout        (),                                                //           (terminated)
		.areset             (1'b0),                                            //           (terminated)
		.locked             (),                                                //           (terminated)
		.phasedone          (),                                                //           (terminated)
		.phasecounterselect (4'b0000),                                         //           (terminated)
		.phaseupdown        (1'b0),                                            //           (terminated)
		.phasestep          (1'b0),                                            //           (terminated)
		.scanclk            (1'b0),                                            //           (terminated)
		.scanclkena         (1'b0),                                            //           (terminated)
		.scandata           (1'b0),                                            //           (terminated)
		.configupdate       (1'b0)                                             //           (terminated)
	);

	lab9_soc_mm_interconnect_0 mm_interconnect_0 (
		.CLK_clk_clk                                (clk_clk),                                                      //                           CLK_clk.clk
		.SDRAM_PLL_c0_clk                           (sdram_pll_c0_clk),                                             //                      SDRAM_PLL_c0.clk
		.NIOS2_reset_reset_bridge_in_reset_reset    (rst_controller_reset_out_reset),                               // NIOS2_reset_reset_bridge_in_reset.reset
		.SDRAM_reset_reset_bridge_in_reset_reset    (rst_controller_001_reset_out_reset),                           // SDRAM_reset_reset_bridge_in_reset.reset
		.NIOS2_data_master_address                  (nios2_data_master_address),                                    //                 NIOS2_data_master.address
		.NIOS2_data_master_waitrequest              (nios2_data_master_waitrequest),                                //                                  .waitrequest
		.NIOS2_data_master_byteenable               (nios2_data_master_byteenable),                                 //                                  .byteenable
		.NIOS2_data_master_read                     (nios2_data_master_read),                                       //                                  .read
		.NIOS2_data_master_readdata                 (nios2_data_master_readdata),                                   //                                  .readdata
		.NIOS2_data_master_write                    (nios2_data_master_write),                                      //                                  .write
		.NIOS2_data_master_writedata                (nios2_data_master_writedata),                                  //                                  .writedata
		.NIOS2_data_master_debugaccess              (nios2_data_master_debugaccess),                                //                                  .debugaccess
		.NIOS2_instruction_master_address           (nios2_instruction_master_address),                             //          NIOS2_instruction_master.address
		.NIOS2_instruction_master_waitrequest       (nios2_instruction_master_waitrequest),                         //                                  .waitrequest
		.NIOS2_instruction_master_read              (nios2_instruction_master_read),                                //                                  .read
		.NIOS2_instruction_master_readdata          (nios2_instruction_master_readdata),                            //                                  .readdata
		.AES_Decryption_Core_0_AES_Slave_address    (mm_interconnect_0_aes_decryption_core_0_aes_slave_address),    //   AES_Decryption_Core_0_AES_Slave.address
		.AES_Decryption_Core_0_AES_Slave_write      (mm_interconnect_0_aes_decryption_core_0_aes_slave_write),      //                                  .write
		.AES_Decryption_Core_0_AES_Slave_read       (mm_interconnect_0_aes_decryption_core_0_aes_slave_read),       //                                  .read
		.AES_Decryption_Core_0_AES_Slave_readdata   (mm_interconnect_0_aes_decryption_core_0_aes_slave_readdata),   //                                  .readdata
		.AES_Decryption_Core_0_AES_Slave_writedata  (mm_interconnect_0_aes_decryption_core_0_aes_slave_writedata),  //                                  .writedata
		.AES_Decryption_Core_0_AES_Slave_byteenable (mm_interconnect_0_aes_decryption_core_0_aes_slave_byteenable), //                                  .byteenable
		.AES_Decryption_Core_0_AES_Slave_chipselect (mm_interconnect_0_aes_decryption_core_0_aes_slave_chipselect), //                                  .chipselect
		.JTAG_UART_avalon_jtag_slave_address        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),        //       JTAG_UART_avalon_jtag_slave.address
		.JTAG_UART_avalon_jtag_slave_write          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),          //                                  .write
		.JTAG_UART_avalon_jtag_slave_read           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),           //                                  .read
		.JTAG_UART_avalon_jtag_slave_readdata       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),       //                                  .readdata
		.JTAG_UART_avalon_jtag_slave_writedata      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),      //                                  .writedata
		.JTAG_UART_avalon_jtag_slave_waitrequest    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),    //                                  .waitrequest
		.JTAG_UART_avalon_jtag_slave_chipselect     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),     //                                  .chipselect
		.NIOS2_debug_mem_slave_address              (mm_interconnect_0_nios2_debug_mem_slave_address),              //             NIOS2_debug_mem_slave.address
		.NIOS2_debug_mem_slave_write                (mm_interconnect_0_nios2_debug_mem_slave_write),                //                                  .write
		.NIOS2_debug_mem_slave_read                 (mm_interconnect_0_nios2_debug_mem_slave_read),                 //                                  .read
		.NIOS2_debug_mem_slave_readdata             (mm_interconnect_0_nios2_debug_mem_slave_readdata),             //                                  .readdata
		.NIOS2_debug_mem_slave_writedata            (mm_interconnect_0_nios2_debug_mem_slave_writedata),            //                                  .writedata
		.NIOS2_debug_mem_slave_byteenable           (mm_interconnect_0_nios2_debug_mem_slave_byteenable),           //                                  .byteenable
		.NIOS2_debug_mem_slave_waitrequest          (mm_interconnect_0_nios2_debug_mem_slave_waitrequest),          //                                  .waitrequest
		.NIOS2_debug_mem_slave_debugaccess          (mm_interconnect_0_nios2_debug_mem_slave_debugaccess),          //                                  .debugaccess
		.NIOS2_SYSID_control_slave_address          (mm_interconnect_0_nios2_sysid_control_slave_address),          //         NIOS2_SYSID_control_slave.address
		.NIOS2_SYSID_control_slave_readdata         (mm_interconnect_0_nios2_sysid_control_slave_readdata),         //                                  .readdata
		.ONCHIP_MEMORY_s1_address                   (mm_interconnect_0_onchip_memory_s1_address),                   //                  ONCHIP_MEMORY_s1.address
		.ONCHIP_MEMORY_s1_write                     (mm_interconnect_0_onchip_memory_s1_write),                     //                                  .write
		.ONCHIP_MEMORY_s1_readdata                  (mm_interconnect_0_onchip_memory_s1_readdata),                  //                                  .readdata
		.ONCHIP_MEMORY_s1_writedata                 (mm_interconnect_0_onchip_memory_s1_writedata),                 //                                  .writedata
		.ONCHIP_MEMORY_s1_byteenable                (mm_interconnect_0_onchip_memory_s1_byteenable),                //                                  .byteenable
		.ONCHIP_MEMORY_s1_chipselect                (mm_interconnect_0_onchip_memory_s1_chipselect),                //                                  .chipselect
		.ONCHIP_MEMORY_s1_clken                     (mm_interconnect_0_onchip_memory_s1_clken),                     //                                  .clken
		.SDRAM_s1_address                           (mm_interconnect_0_sdram_s1_address),                           //                          SDRAM_s1.address
		.SDRAM_s1_write                             (mm_interconnect_0_sdram_s1_write),                             //                                  .write
		.SDRAM_s1_read                              (mm_interconnect_0_sdram_s1_read),                              //                                  .read
		.SDRAM_s1_readdata                          (mm_interconnect_0_sdram_s1_readdata),                          //                                  .readdata
		.SDRAM_s1_writedata                         (mm_interconnect_0_sdram_s1_writedata),                         //                                  .writedata
		.SDRAM_s1_byteenable                        (mm_interconnect_0_sdram_s1_byteenable),                        //                                  .byteenable
		.SDRAM_s1_readdatavalid                     (mm_interconnect_0_sdram_s1_readdatavalid),                     //                                  .readdatavalid
		.SDRAM_s1_waitrequest                       (mm_interconnect_0_sdram_s1_waitrequest),                       //                                  .waitrequest
		.SDRAM_s1_chipselect                        (mm_interconnect_0_sdram_s1_chipselect),                        //                                  .chipselect
		.SDRAM_PLL_pll_slave_address                (mm_interconnect_0_sdram_pll_pll_slave_address),                //               SDRAM_PLL_pll_slave.address
		.SDRAM_PLL_pll_slave_write                  (mm_interconnect_0_sdram_pll_pll_slave_write),                  //                                  .write
		.SDRAM_PLL_pll_slave_read                   (mm_interconnect_0_sdram_pll_pll_slave_read),                   //                                  .read
		.SDRAM_PLL_pll_slave_readdata               (mm_interconnect_0_sdram_pll_pll_slave_readdata),               //                                  .readdata
		.SDRAM_PLL_pll_slave_writedata              (mm_interconnect_0_sdram_pll_pll_slave_writedata)               //                                  .writedata
	);

	lab9_soc_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios2_debug_reset_request_reset),    // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios2_debug_reset_request_reset),    // reset_in1.reset
		.clk            (sdram_pll_c0_clk),                   //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
