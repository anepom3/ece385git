module ShooterSprite (
	input  logic clk,
	input  logic [9:0] in,
	output logic [23:0] out
);

// This module will be synthesized into a RAM
always_ff @ (negedge clk)
	case (in)
  10'h000: out <= 24'hffffff;    10'h080: out <= 24'hffffff;    10'h100: out <= 24'hffffff;    10'h180: out <= 24'hffffff;    10'h200: out <= 24'hffffff;    10'h280: out <= 24'h8a6e47;    10'h300: out <= 24'hffffff;    10'h380: out <= 24'hffffff;
  10'h001: out <= 24'hffffff;    10'h081: out <= 24'hffffff;    10'h101: out <= 24'hffffff;    10'h181: out <= 24'hffffff;    10'h201: out <= 24'hffffff;    10'h281: out <= 24'hffffff;    10'h301: out <= 24'hffffff;    10'h381: out <= 24'hffffff;
  10'h002: out <= 24'hffffff;    10'h082: out <= 24'hffffff;    10'h102: out <= 24'hffffff;    10'h182: out <= 24'hffffff;    10'h202: out <= 24'h000000;    10'h282: out <= 24'hffffff;    10'h302: out <= 24'h000000;    10'h382: out <= 24'hffffff;
  10'h003: out <= 24'hffffff;    10'h083: out <= 24'hffffff;    10'h103: out <= 24'hffffff;    10'h183: out <= 24'hffffff;    10'h203: out <= 24'h8a6e47;    10'h283: out <= 24'h000000;    10'h303: out <= 24'h8a6e47;    10'h383: out <= 24'h000000;
  10'h004: out <= 24'hffffff;    10'h084: out <= 24'hffffff;    10'h104: out <= 24'hffffff;    10'h184: out <= 24'h000000;    10'h204: out <= 24'h404f2c;    10'h284: out <= 24'h8a6e47;    10'h304: out <= 24'h404f2c;    10'h384: out <= 24'h8a6e47;
  10'h005: out <= 24'hffffff;    10'h085: out <= 24'hffffff;    10'h105: out <= 24'hffffff;    10'h185: out <= 24'h8a6e47;    10'h205: out <= 24'h8a6e47;    10'h285: out <= 24'h404f2c;    10'h305: out <= 24'h8a6e47;    10'h385: out <= 24'h8a6e47;
  10'h006: out <= 24'hffffff;    10'h086: out <= 24'hffffff;    10'h106: out <= 24'hffffff;    10'h186: out <= 24'h8a6e47;    10'h206: out <= 24'h8a6e47;    10'h286: out <= 24'h404f2c;    10'h306: out <= 24'h8a6e47;    10'h386: out <= 24'h8a6e47;
  10'h007: out <= 24'hffffff;    10'h087: out <= 24'hffffff;    10'h107: out <= 24'h000000;    10'h187: out <= 24'h8a6e47;    10'h207: out <= 24'h8a6e47;    10'h287: out <= 24'h8a6e47;    10'h307: out <= 24'h8a6e47;    10'h387: out <= 24'h8a6e47;
  10'h008: out <= 24'hffffff;    10'h088: out <= 24'hffffff;    10'h108: out <= 24'h000000;    10'h188: out <= 24'h8a6e47;    10'h208: out <= 24'h8a6e47;    10'h288: out <= 24'h8a6e47;    10'h308: out <= 24'h000000;    10'h388: out <= 24'h8a6e47;
  10'h009: out <= 24'hffffff;    10'h089: out <= 24'hffffff;    10'h109: out <= 24'h404f2c;    10'h189: out <= 24'h8a6e47;    10'h209: out <= 24'h000000;    10'h289: out <= 24'h000000;    10'h309: out <= 24'hffffff;    10'h389: out <= 24'h8a6e47;
  10'h00a: out <= 24'hffffff;    10'h08a: out <= 24'hffffff;    10'h10a: out <= 24'h8a6e47;    10'h18a: out <= 24'h000000;    10'h20a: out <= 24'hffffff;    10'h28a: out <= 24'hffffff;    10'h30a: out <= 24'h000000;    10'h38a: out <= 24'h000000;
  10'h00b: out <= 24'hffffff;    10'h08b: out <= 24'hffffff;    10'h10b: out <= 24'h8a6e47;    10'h18b: out <= 24'h000000;    10'h20b: out <= 24'hffffff;    10'h28b: out <= 24'hffffff;    10'h30b: out <= 24'h8a6e47;    10'h38b: out <= 24'h886028;
  10'h00c: out <= 24'hffffff;    10'h08c: out <= 24'h000000;    10'h10c: out <= 24'h8a6e47;    10'h18c: out <= 24'hffffff;    10'h20c: out <= 24'hffffff;    10'h28c: out <= 24'hffffff;    10'h30c: out <= 24'h000000;    10'h38c: out <= 24'h886028;
  10'h00d: out <= 24'hffffff;    10'h08d: out <= 24'h6c4a1b;    10'h10d: out <= 24'h8a6e47;    10'h18d: out <= 24'hffffff;    10'h20d: out <= 24'hffffff;    10'h28d: out <= 24'h000000;    10'h30d: out <= 24'hffc18f;    10'h38d: out <= 24'h886028;
  10'h00e: out <= 24'hffffff;    10'h08e: out <= 24'h6c4a1b;    10'h10e: out <= 24'h000000;    10'h18e: out <= 24'hffffff;    10'h20e: out <= 24'hffffff;    10'h28e: out <= 24'h8a6e47;    10'h30e: out <= 24'hffc18f;    10'h38e: out <= 24'h886028;
  10'h00f: out <= 24'hffffff;    10'h08f: out <= 24'h000000;    10'h10f: out <= 24'hffffff;    10'h18f: out <= 24'hffffff;    10'h20f: out <= 24'hffffff;    10'h28f: out <= 24'h404f2c;    10'h30f: out <= 24'hffc18f;    10'h38f: out <= 24'h886028;
  10'h010: out <= 24'h000000;    10'h090: out <= 24'h000000;    10'h110: out <= 24'hffffff;    10'h190: out <= 24'hffffff;    10'h210: out <= 24'hffffff;    10'h290: out <= 24'h404f2c;    10'h310: out <= 24'hffc18f;    10'h390: out <= 24'h886028;
  10'h011: out <= 24'hffffff;    10'h091: out <= 24'h000000;    10'h111: out <= 24'hffffff;    10'h191: out <= 24'hffffff;    10'h211: out <= 24'hffffff;    10'h291: out <= 24'h8a6e47;    10'h311: out <= 24'hffc18f;    10'h391: out <= 24'h886028;
  10'h012: out <= 24'hffffff;    10'h092: out <= 24'h6c4a1b;    10'h112: out <= 24'h000000;    10'h192: out <= 24'hffffff;    10'h212: out <= 24'hffffff;    10'h292: out <= 24'h8a6e47;    10'h312: out <= 24'hffc18f;    10'h392: out <= 24'h886028;
  10'h013: out <= 24'hffffff;    10'h093: out <= 24'h6c4a1b;    10'h113: out <= 24'h8a6e47;    10'h193: out <= 24'hffffff;    10'h213: out <= 24'hffffff;    10'h293: out <= 24'h404f2c;    10'h313: out <= 24'h000000;    10'h393: out <= 24'h886028;
  10'h014: out <= 24'hffffff;    10'h094: out <= 24'h000000;    10'h114: out <= 24'h8a6e47;    10'h194: out <= 24'hffffff;    10'h214: out <= 24'hffffff;    10'h294: out <= 24'h000000;    10'h314: out <= 24'h8a6e47;    10'h394: out <= 24'h886028;
  10'h015: out <= 24'hffffff;    10'h095: out <= 24'hffffff;    10'h115: out <= 24'h8a6e47;    10'h195: out <= 24'h000000;    10'h215: out <= 24'hffffff;    10'h295: out <= 24'hffffff;    10'h315: out <= 24'h000000;    10'h395: out <= 24'h000000;
  10'h016: out <= 24'hffffff;    10'h096: out <= 24'hffffff;    10'h116: out <= 24'h8a6e47;    10'h196: out <= 24'h404f2c;    10'h216: out <= 24'hffffff;    10'h296: out <= 24'hffffff;    10'h316: out <= 24'hffffff;    10'h396: out <= 24'h8a6e47;
  10'h017: out <= 24'hffffff;    10'h097: out <= 24'hffffff;    10'h117: out <= 24'h8a6e47;    10'h197: out <= 24'h8a6e47;    10'h217: out <= 24'h000000;    10'h297: out <= 24'hffffff;    10'h317: out <= 24'h000000;    10'h397: out <= 24'h8a6e47;
  10'h018: out <= 24'hffffff;    10'h098: out <= 24'hffffff;    10'h118: out <= 24'h000000;    10'h198: out <= 24'h8a6e47;    10'h218: out <= 24'h404f2c;    10'h298: out <= 24'h000000;    10'h318: out <= 24'h8a6e47;    10'h398: out <= 24'h8a6e47;
  10'h019: out <= 24'hffffff;    10'h099: out <= 24'hffffff;    10'h119: out <= 24'h000000;    10'h199: out <= 24'h8a6e47;    10'h219: out <= 24'h8a6e47;    10'h299: out <= 24'h8a6e47;    10'h319: out <= 24'h8a6e47;    10'h399: out <= 24'h8a6e47;
  10'h01a: out <= 24'hffffff;    10'h09a: out <= 24'hffffff;    10'h11a: out <= 24'hffffff;    10'h19a: out <= 24'h8a6e47;    10'h21a: out <= 24'h8a6e47;    10'h29a: out <= 24'h8a6e47;    10'h31a: out <= 24'h8a6e47;    10'h39a: out <= 24'h8a6e47;
  10'h01b: out <= 24'hffffff;    10'h09b: out <= 24'hffffff;    10'h11b: out <= 24'hffffff;    10'h19b: out <= 24'h000000;    10'h21b: out <= 24'h8a6e47;    10'h29b: out <= 24'h8a6e47;    10'h31b: out <= 24'h8a6e47;    10'h39b: out <= 24'h8a6e47;
  10'h01c: out <= 24'hffffff;    10'h09c: out <= 24'hffffff;    10'h11c: out <= 24'hffffff;    10'h19c: out <= 24'h000000;    10'h21c: out <= 24'h8a6e47;    10'h29c: out <= 24'h404f2c;    10'h31c: out <= 24'h8a6e47;    10'h39c: out <= 24'h000000;
  10'h01d: out <= 24'hffffff;    10'h09d: out <= 24'hffffff;    10'h11d: out <= 24'hffffff;    10'h19d: out <= 24'hffffff;    10'h21d: out <= 24'h000000;    10'h29d: out <= 24'h000000;    10'h31d: out <= 24'h000000;    10'h39d: out <= 24'hffffff;
  10'h01e: out <= 24'hffffff;    10'h09e: out <= 24'hffffff;    10'h11e: out <= 24'hffffff;    10'h19e: out <= 24'hffffff;    10'h21e: out <= 24'hffffff;    10'h29e: out <= 24'hffffff;    10'h31e: out <= 24'hffffff;    10'h39e: out <= 24'hffffff;
  10'h01f: out <= 24'hffffff;    10'h09f: out <= 24'hffffff;    10'h11f: out <= 24'hffffff;    10'h19f: out <= 24'hffffff;    10'h21f: out <= 24'hffffff;    10'h29f: out <= 24'hffffff;    10'h31f: out <= 24'hffffff;    10'h39f: out <= 24'hffffff;
  10'h020: out <= 24'hffffff;    10'h0a0: out <= 24'hffffff;    10'h120: out <= 24'hffffff;    10'h1a0: out <= 24'hffffff;    10'h220: out <= 24'hffffff;    10'h2a0: out <= 24'hffffff;    10'h320: out <= 24'hffffff;    10'h3a0: out <= 24'hffffff;
  10'h021: out <= 24'hffffff;    10'h0a1: out <= 24'hffffff;    10'h121: out <= 24'hffffff;    10'h1a1: out <= 24'hffffff;    10'h221: out <= 24'hffffff;    10'h2a1: out <= 24'hffffff;    10'h321: out <= 24'hffffff;    10'h3a1: out <= 24'hffffff;
  10'h022: out <= 24'hffffff;    10'h0a2: out <= 24'hffffff;    10'h122: out <= 24'hffffff;    10'h1a2: out <= 24'hffffff;    10'h222: out <= 24'h000000;    10'h2a2: out <= 24'h000000;    10'h322: out <= 24'h000000;    10'h3a2: out <= 24'hffffff;
  10'h023: out <= 24'hffffff;    10'h0a3: out <= 24'hffffff;    10'h123: out <= 24'hffffff;    10'h1a3: out <= 24'h000000;    10'h223: out <= 24'h404f2c;    10'h2a3: out <= 24'h8a6e47;    10'h323: out <= 24'h8a6e47;    10'h3a3: out <= 24'hffffff;
  10'h024: out <= 24'hffffff;    10'h0a4: out <= 24'hffffff;    10'h124: out <= 24'hffffff;    10'h1a4: out <= 24'h404f2c;    10'h224: out <= 24'h404f2c;    10'h2a4: out <= 24'h8a6e47;    10'h324: out <= 24'h8a6e47;    10'h3a4: out <= 24'h000000;
  10'h025: out <= 24'hffffff;    10'h0a5: out <= 24'hffffff;    10'h125: out <= 24'hffffff;    10'h1a5: out <= 24'h404f2c;    10'h225: out <= 24'h8a6e47;    10'h2a5: out <= 24'h8a6e47;    10'h325: out <= 24'h8a6e47;    10'h3a5: out <= 24'h8a6e47;
  10'h026: out <= 24'hffffff;    10'h0a6: out <= 24'hffffff;    10'h126: out <= 24'h000000;    10'h1a6: out <= 24'h8a6e47;    10'h226: out <= 24'h8a6e47;    10'h2a6: out <= 24'h8a6e47;    10'h326: out <= 24'h8a6e47;    10'h3a6: out <= 24'h8a6e47;
  10'h027: out <= 24'hffffff;    10'h0a7: out <= 24'hffffff;    10'h127: out <= 24'h000000;    10'h1a7: out <= 24'h8a6e47;    10'h227: out <= 24'h404f2c;    10'h2a7: out <= 24'h8a6e47;    10'h327: out <= 24'h8a6e47;    10'h3a7: out <= 24'h8a6e47;
  10'h028: out <= 24'hffffff;    10'h0a8: out <= 24'hffffff;    10'h128: out <= 24'h8a6e47;    10'h1a8: out <= 24'h8a6e47;    10'h228: out <= 24'h000000;    10'h2a8: out <= 24'h000000;    10'h328: out <= 24'h000000;    10'h3a8: out <= 24'h404f2c;
  10'h029: out <= 24'hffffff;    10'h0a9: out <= 24'hffffff;    10'h129: out <= 24'h404f2c;    10'h1a9: out <= 24'h404f2c;    10'h229: out <= 24'hffffff;    10'h2a9: out <= 24'hffffff;    10'h329: out <= 24'hffffff;    10'h3a9: out <= 24'h8a6e47;
  10'h02a: out <= 24'hffffff;    10'h0aa: out <= 24'h000000;    10'h12a: out <= 24'h8a6e47;    10'h1aa: out <= 24'h000000;    10'h22a: out <= 24'hffffff;    10'h2aa: out <= 24'hffffff;    10'h32a: out <= 24'h000000;    10'h3aa: out <= 24'h8a6e47;
  10'h02b: out <= 24'hffffff;    10'h0ab: out <= 24'h000000;    10'h12b: out <= 24'h8a6e47;    10'h1ab: out <= 24'hffffff;    10'h22b: out <= 24'hffffff;    10'h2ab: out <= 24'h000000;    10'h32b: out <= 24'h000000;    10'h3ab: out <= 24'h000000;
  10'h02c: out <= 24'hffffff;    10'h0ac: out <= 24'h000000;    10'h12c: out <= 24'h8a6e47;    10'h1ac: out <= 24'hffffff;    10'h22c: out <= 24'hffffff;    10'h2ac: out <= 24'h8a6e47;    10'h32c: out <= 24'hffc18f;    10'h3ac: out <= 24'h886028;
  10'h02d: out <= 24'hffffff;    10'h0ad: out <= 24'h6c4a1b;    10'h12d: out <= 24'h000000;    10'h1ad: out <= 24'hffffff;    10'h22d: out <= 24'hffffff;    10'h2ad: out <= 24'h8a6e47;    10'h32d: out <= 24'hffc18f;    10'h3ad: out <= 24'h886028;
  10'h02e: out <= 24'hffffff;    10'h0ae: out <= 24'h6c4a1b;    10'h12e: out <= 24'h000000;    10'h1ae: out <= 24'hffffff;    10'h22e: out <= 24'hffffff;    10'h2ae: out <= 24'h8a6e47;    10'h32e: out <= 24'h000000;    10'h3ae: out <= 24'h886028;
  10'h02f: out <= 24'h000000;    10'h0af: out <= 24'h000000;    10'h12f: out <= 24'hffffff;    10'h1af: out <= 24'hffffff;    10'h22f: out <= 24'hffffff;    10'h2af: out <= 24'h8a6e47;    10'h32f: out <= 24'hffc18f;    10'h3af: out <= 24'h886028;
  10'h030: out <= 24'h000000;    10'h0b0: out <= 24'h000000;    10'h130: out <= 24'hffffff;    10'h1b0: out <= 24'hffffff;    10'h230: out <= 24'hffffff;    10'h2b0: out <= 24'h8a6e47;    10'h330: out <= 24'hffc18f;    10'h3b0: out <= 24'h886028;
  10'h031: out <= 24'h000000;    10'h0b1: out <= 24'h000000;    10'h131: out <= 24'hffffff;    10'h1b1: out <= 24'hffffff;    10'h231: out <= 24'hffffff;    10'h2b1: out <= 24'h8a6e47;    10'h331: out <= 24'h000000;    10'h3b1: out <= 24'h886028;
  10'h032: out <= 24'hffffff;    10'h0b2: out <= 24'h6c4a1b;    10'h132: out <= 24'h000000;    10'h1b2: out <= 24'hffffff;    10'h232: out <= 24'hffffff;    10'h2b2: out <= 24'h8a6e47;    10'h332: out <= 24'hffc18f;    10'h3b2: out <= 24'h886028;
  10'h033: out <= 24'hffffff;    10'h0b3: out <= 24'h6c4a1b;    10'h133: out <= 24'h000000;    10'h1b3: out <= 24'hffffff;    10'h233: out <= 24'hffffff;    10'h2b3: out <= 24'h404f2c;    10'h333: out <= 24'hffc18f;    10'h3b3: out <= 24'h886028;
  10'h034: out <= 24'hffffff;    10'h0b4: out <= 24'h000000;    10'h134: out <= 24'h8a6e47;    10'h1b4: out <= 24'hffffff;    10'h234: out <= 24'hffffff;    10'h2b4: out <= 24'h000000;    10'h334: out <= 24'h000000;    10'h3b4: out <= 24'h000000;
  10'h035: out <= 24'hffffff;    10'h0b5: out <= 24'h000000;    10'h135: out <= 24'h8a6e47;    10'h1b5: out <= 24'h000000;    10'h235: out <= 24'hffffff;    10'h2b5: out <= 24'hffffff;    10'h335: out <= 24'h000000;    10'h3b5: out <= 24'h8a6e47;
  10'h036: out <= 24'hffffff;    10'h0b6: out <= 24'h000000;    10'h136: out <= 24'h8a6e47;    10'h1b6: out <= 24'h000000;    10'h236: out <= 24'hffffff;    10'h2b6: out <= 24'hffffff;    10'h336: out <= 24'hffffff;    10'h3b6: out <= 24'h8a6e47;
  10'h037: out <= 24'hffffff;    10'h0b7: out <= 24'hffffff;    10'h137: out <= 24'h8a6e47;    10'h1b7: out <= 24'h404f2c;    10'h237: out <= 24'h000000;    10'h2b7: out <= 24'h000000;    10'h337: out <= 24'h000000;    10'h3b7: out <= 24'h8a6e47;
  10'h038: out <= 24'hffffff;    10'h0b8: out <= 24'hffffff;    10'h138: out <= 24'h8a6e47;    10'h1b8: out <= 24'h8a6e47;    10'h238: out <= 24'h404f2c;    10'h2b8: out <= 24'h8a6e47;    10'h338: out <= 24'h8a6e47;    10'h3b8: out <= 24'h8a6e47;
  10'h039: out <= 24'hffffff;    10'h0b9: out <= 24'hffffff;    10'h139: out <= 24'h000000;    10'h1b9: out <= 24'h8a6e47;    10'h239: out <= 24'h8a6e47;    10'h2b9: out <= 24'h8a6e47;    10'h339: out <= 24'h8a6e47;    10'h3b9: out <= 24'h8a6e47;
  10'h03a: out <= 24'hffffff;    10'h0ba: out <= 24'hffffff;    10'h13a: out <= 24'h000000;    10'h1ba: out <= 24'h8a6e47;    10'h23a: out <= 24'h8a6e47;    10'h2ba: out <= 24'h8a6e47;    10'h33a: out <= 24'h8a6e47;    10'h3ba: out <= 24'h8a6e47;
  10'h03b: out <= 24'hffffff;    10'h0bb: out <= 24'hffffff;    10'h13b: out <= 24'hffffff;    10'h1bb: out <= 24'h404f2c;    10'h23b: out <= 24'h404f2c;    10'h2bb: out <= 24'h8a6e47;    10'h33b: out <= 24'h8a6e47;    10'h3bb: out <= 24'h000000;
  10'h03c: out <= 24'hffffff;    10'h0bc: out <= 24'hffffff;    10'h13c: out <= 24'hffffff;    10'h1bc: out <= 24'h000000;    10'h23c: out <= 24'h404f2c;    10'h2bc: out <= 24'h8a6e47;    10'h33c: out <= 24'h8a6e47;    10'h3bc: out <= 24'hffffff;
  10'h03d: out <= 24'hffffff;    10'h0bd: out <= 24'hffffff;    10'h13d: out <= 24'hffffff;    10'h1bd: out <= 24'hffffff;    10'h23d: out <= 24'h000000;    10'h2bd: out <= 24'h000000;    10'h33d: out <= 24'h000000;    10'h3bd: out <= 24'hffffff;
  10'h03e: out <= 24'hffffff;    10'h0be: out <= 24'hffffff;    10'h13e: out <= 24'hffffff;    10'h1be: out <= 24'hffffff;    10'h23e: out <= 24'hffffff;    10'h2be: out <= 24'hffffff;    10'h33e: out <= 24'hffffff;    10'h3be: out <= 24'hffffff;
  10'h03f: out <= 24'hffffff;    10'h0bf: out <= 24'hffffff;    10'h13f: out <= 24'hffffff;    10'h1bf: out <= 24'hffffff;    10'h23f: out <= 24'hffffff;    10'h2bf: out <= 24'hffffff;    10'h33f: out <= 24'hffffff;    10'h3bf: out <= 24'hffffff;
  10'h040: out <= 24'hffffff;    10'h0c0: out <= 24'hffffff;    10'h140: out <= 24'hffffff;    10'h1c0: out <= 24'hffffff;    10'h240: out <= 24'hffffff;    10'h2c0: out <= 24'hffffff;    10'h340: out <= 24'hffffff;    10'h3c0: out <= 24'hffffff;
  10'h041: out <= 24'hffffff;    10'h0c1: out <= 24'hffffff;    10'h141: out <= 24'hffffff;    10'h1c1: out <= 24'hffffff;    10'h241: out <= 24'hffffff;    10'h2c1: out <= 24'hffffff;    10'h341: out <= 24'hffffff;    10'h3c1: out <= 24'hffffff;
  10'h042: out <= 24'hffffff;    10'h0c2: out <= 24'hffffff;    10'h142: out <= 24'hffffff;    10'h1c2: out <= 24'hffffff;    10'h242: out <= 24'h000000;    10'h2c2: out <= 24'h000000;    10'h342: out <= 24'h000000;    10'h3c2: out <= 24'hffffff;
  10'h043: out <= 24'hffffff;    10'h0c3: out <= 24'hffffff;    10'h143: out <= 24'hffffff;    10'h1c3: out <= 24'h000000;    10'h243: out <= 24'h8a6e47;    10'h2c3: out <= 24'h8a6e47;    10'h343: out <= 24'h8a6e47;    10'h3c3: out <= 24'hffffff;
  10'h044: out <= 24'hffffff;    10'h0c4: out <= 24'hffffff;    10'h144: out <= 24'hffffff;    10'h1c4: out <= 24'h8a6e47;    10'h244: out <= 24'h8a6e47;    10'h2c4: out <= 24'h8a6e47;    10'h344: out <= 24'h8a6e47;    10'h3c4: out <= 24'hffffff;
  10'h045: out <= 24'hffffff;    10'h0c5: out <= 24'hffffff;    10'h145: out <= 24'h000000;    10'h1c5: out <= 24'h8a6e47;    10'h245: out <= 24'h8a6e47;    10'h2c5: out <= 24'h8a6e47;    10'h345: out <= 24'h8a6e47;    10'h3c5: out <= 24'h000000;
  10'h046: out <= 24'hffffff;    10'h0c6: out <= 24'hffffff;    10'h146: out <= 24'h000000;    10'h1c6: out <= 24'h8a6e47;    10'h246: out <= 24'h8a6e47;    10'h2c6: out <= 24'h8a6e47;    10'h346: out <= 24'h8a6e47;    10'h3c6: out <= 24'h8a6e47;
  10'h047: out <= 24'hffffff;    10'h0c7: out <= 24'hffffff;    10'h147: out <= 24'h8a6e47;    10'h1c7: out <= 24'h8a6e47;    10'h247: out <= 24'h404f2c;    10'h2c7: out <= 24'h8a6e47;    10'h347: out <= 24'h8a6e47;    10'h3c7: out <= 24'h8a6e47;
  10'h048: out <= 24'hffffff;    10'h0c8: out <= 24'hffffff;    10'h148: out <= 24'h8a6e47;    10'h1c8: out <= 24'h404f2c;    10'h248: out <= 24'h000000;    10'h2c8: out <= 24'h000000;    10'h348: out <= 24'h404f2c;    10'h3c8: out <= 24'h404f2c;
  10'h049: out <= 24'hffffff;    10'h0c9: out <= 24'h000000;    10'h149: out <= 24'h8a6e47;    10'h1c9: out <= 24'h000000;    10'h249: out <= 24'hffffff;    10'h2c9: out <= 24'hffffff;    10'h349: out <= 24'h000000;    10'h3c9: out <= 24'h8a6e47;
  10'h04a: out <= 24'hffffff;    10'h0ca: out <= 24'h000000;    10'h14a: out <= 24'h8a6e47;    10'h1ca: out <= 24'h000000;    10'h24a: out <= 24'hffffff;    10'h2ca: out <= 24'h000000;    10'h34a: out <= 24'h000000;    10'h3ca: out <= 24'h8a6e47;
  10'h04b: out <= 24'hffffff;    10'h0cb: out <= 24'h8a6e47;    10'h14b: out <= 24'h8a6e47;    10'h1cb: out <= 24'hffffff;    10'h24b: out <= 24'hffffff;    10'h2cb: out <= 24'h404f2c;    10'h34b: out <= 24'hffc18f;    10'h3cb: out <= 24'h8a6e47;
  10'h04c: out <= 24'hffffff;    10'h0cc: out <= 24'h000000;    10'h14c: out <= 24'h000000;    10'h1cc: out <= 24'hffffff;    10'h24c: out <= 24'hffffff;    10'h2cc: out <= 24'h404f2c;    10'h34c: out <= 24'hffc18f;    10'h3cc: out <= 24'h000000;
  10'h04d: out <= 24'hffffff;    10'h0cd: out <= 24'h6c4a1b;    10'h14d: out <= 24'h000000;    10'h1cd: out <= 24'hffffff;    10'h24d: out <= 24'hffffff;    10'h2cd: out <= 24'h8a6e47;    10'h34d: out <= 24'hffc18f;    10'h3cd: out <= 24'h886028;
  10'h04e: out <= 24'hffffff;    10'h0ce: out <= 24'h6c4a1b;    10'h14e: out <= 24'hffffff;    10'h1ce: out <= 24'hffffff;    10'h24e: out <= 24'hffffff;    10'h2ce: out <= 24'h8a6e47;    10'h34e: out <= 24'hffc18f;    10'h3ce: out <= 24'h886028;
  10'h04f: out <= 24'h000000;    10'h0cf: out <= 24'h6c4a1b;    10'h14f: out <= 24'hffffff;    10'h1cf: out <= 24'hffffff;    10'h24f: out <= 24'hffffff;    10'h2cf: out <= 24'h000000;    10'h34f: out <= 24'hffc18f;    10'h3cf: out <= 24'h886028;
  10'h050: out <= 24'h000000;    10'h0d0: out <= 24'h000000;    10'h150: out <= 24'hffffff;    10'h1d0: out <= 24'hffffff;    10'h250: out <= 24'hffffff;    10'h2d0: out <= 24'h000000;    10'h350: out <= 24'hffc18f;    10'h3d0: out <= 24'h886028;
  10'h051: out <= 24'h000000;    10'h0d1: out <= 24'h6c4a1b;    10'h151: out <= 24'hffffff;    10'h1d1: out <= 24'hffffff;    10'h251: out <= 24'hffffff;    10'h2d1: out <= 24'h8a6e47;    10'h351: out <= 24'hffc18f;    10'h3d1: out <= 24'h886028;
  10'h052: out <= 24'hffffff;    10'h0d2: out <= 24'h6c4a1b;    10'h152: out <= 24'hffffff;    10'h1d2: out <= 24'hffffff;    10'h252: out <= 24'hffffff;    10'h2d2: out <= 24'h8a6e47;    10'h352: out <= 24'hffc18f;    10'h3d2: out <= 24'h886028;
  10'h053: out <= 24'hffffff;    10'h0d3: out <= 24'h6c4a1b;    10'h153: out <= 24'hffffff;    10'h1d3: out <= 24'hffffff;    10'h253: out <= 24'hffffff;    10'h2d3: out <= 24'h8a6e47;    10'h353: out <= 24'hffc18f;    10'h3d3: out <= 24'h000000;
  10'h054: out <= 24'hffffff;    10'h0d4: out <= 24'h000000;    10'h154: out <= 24'h000000;    10'h1d4: out <= 24'hffffff;    10'h254: out <= 24'hffffff;    10'h2d4: out <= 24'h8a6e47;    10'h354: out <= 24'hffc18f;    10'h3d4: out <= 24'h8a6e47;
  10'h055: out <= 24'hffffff;    10'h0d5: out <= 24'h8a6e47;    10'h155: out <= 24'h8a6e47;    10'h1d5: out <= 24'hffffff;    10'h255: out <= 24'hffffff;    10'h2d5: out <= 24'h000000;    10'h355: out <= 24'h000000;    10'h3d5: out <= 24'h8a6e47;
  10'h056: out <= 24'hffffff;    10'h0d6: out <= 24'h000000;    10'h156: out <= 24'h8a6e47;    10'h1d6: out <= 24'h000000;    10'h256: out <= 24'hffffff;    10'h2d6: out <= 24'hffffff;    10'h356: out <= 24'h000000;    10'h3d6: out <= 24'h8a6e47;
  10'h057: out <= 24'hffffff;    10'h0d7: out <= 24'h000000;    10'h157: out <= 24'h8a6e47;    10'h1d7: out <= 24'h8a6e47;    10'h257: out <= 24'h000000;    10'h2d7: out <= 24'h000000;    10'h357: out <= 24'h404f2c;    10'h3d7: out <= 24'h8a6e47;
  10'h058: out <= 24'hffffff;    10'h0d8: out <= 24'hffffff;    10'h158: out <= 24'h404f2c;    10'h1d8: out <= 24'h8a6e47;    10'h258: out <= 24'h404f2c;    10'h2d8: out <= 24'h8a6e47;    10'h358: out <= 24'h8a6e47;    10'h3d8: out <= 24'h404f2c;
  10'h059: out <= 24'hffffff;    10'h0d9: out <= 24'hffffff;    10'h159: out <= 24'h404f2c;    10'h1d9: out <= 24'h8a6e47;    10'h259: out <= 24'h8a6e47;    10'h2d9: out <= 24'h404f2c;    10'h359: out <= 24'h8a6e47;    10'h3d9: out <= 24'h404f2c;
  10'h05a: out <= 24'hffffff;    10'h0da: out <= 24'hffffff;    10'h15a: out <= 24'h000000;    10'h1da: out <= 24'h404f2c;    10'h25a: out <= 24'h8a6e47;    10'h2da: out <= 24'h404f2c;    10'h35a: out <= 24'h8a6e47;    10'h3da: out <= 24'h000000;
  10'h05b: out <= 24'hffffff;    10'h0db: out <= 24'hffffff;    10'h15b: out <= 24'h000000;    10'h1db: out <= 24'h8a6e47;    10'h25b: out <= 24'h404f2c;    10'h2db: out <= 24'h8a6e47;    10'h35b: out <= 24'h8a6e47;    10'h3db: out <= 24'hffffff;
  10'h05c: out <= 24'hffffff;    10'h0dc: out <= 24'hffffff;    10'h15c: out <= 24'hffffff;    10'h1dc: out <= 24'h000000;    10'h25c: out <= 24'h8a6e47;    10'h2dc: out <= 24'h8a6e47;    10'h35c: out <= 24'h8a6e47;    10'h3dc: out <= 24'hffffff;
  10'h05d: out <= 24'hffffff;    10'h0dd: out <= 24'hffffff;    10'h15d: out <= 24'hffffff;    10'h1dd: out <= 24'hffffff;    10'h25d: out <= 24'h000000;    10'h2dd: out <= 24'h000000;    10'h35d: out <= 24'h000000;    10'h3dd: out <= 24'hffffff;
  10'h05e: out <= 24'hffffff;    10'h0de: out <= 24'hffffff;    10'h15e: out <= 24'hffffff;    10'h1de: out <= 24'hffffff;    10'h25e: out <= 24'hffffff;    10'h2de: out <= 24'hffffff;    10'h35e: out <= 24'hffffff;    10'h3de: out <= 24'hffffff;
  10'h05f: out <= 24'hffffff;    10'h0df: out <= 24'hffffff;    10'h15f: out <= 24'hffffff;    10'h1df: out <= 24'hffffff;    10'h25f: out <= 24'hffffff;    10'h2df: out <= 24'hffffff;    10'h35f: out <= 24'hffffff;    10'h3df: out <= 24'hffffff;
  10'h060: out <= 24'hffffff;    10'h0e0: out <= 24'hffffff;    10'h160: out <= 24'hffffff;    10'h1e0: out <= 24'hffffff;    10'h260: out <= 24'hffffff;    10'h2e0: out <= 24'hffffff;    10'h360: out <= 24'hffffff;    10'h3e0: out <= 24'hffffff;
  10'h061: out <= 24'hffffff;    10'h0e1: out <= 24'hffffff;    10'h161: out <= 24'hffffff;    10'h1e1: out <= 24'hffffff;    10'h261: out <= 24'hffffff;    10'h2e1: out <= 24'hffffff;    10'h361: out <= 24'hffffff;    10'h3e1: out <= 24'hffffff;
  10'h062: out <= 24'hffffff;    10'h0e2: out <= 24'hffffff;    10'h162: out <= 24'hffffff;    10'h1e2: out <= 24'hffffff;    10'h262: out <= 24'h000000;    10'h2e2: out <= 24'h000000;    10'h362: out <= 24'h000000;    10'h3e2: out <= 24'hffffff;
  10'h063: out <= 24'hffffff;    10'h0e3: out <= 24'hffffff;    10'h163: out <= 24'hffffff;    10'h1e3: out <= 24'h000000;    10'h263: out <= 24'h8a6e47;    10'h2e3: out <= 24'h8a6e47;    10'h363: out <= 24'h8a6e47;    10'h3e3: out <= 24'hffffff;
  10'h064: out <= 24'hffffff;    10'h0e4: out <= 24'hffffff;    10'h164: out <= 24'h000000;    10'h1e4: out <= 24'h8a6e47;    10'h264: out <= 24'h8a6e47;    10'h2e4: out <= 24'h8a6e47;    10'h364: out <= 24'h404f2c;    10'h3e4: out <= 24'hffffff;
  10'h065: out <= 24'hffffff;    10'h0e5: out <= 24'hffffff;    10'h165: out <= 24'h000000;    10'h1e5: out <= 24'h8a6e47;    10'h265: out <= 24'h8a6e47;    10'h2e5: out <= 24'h8a6e47;    10'h365: out <= 24'h8a6e47;    10'h3e5: out <= 24'h000000;
  10'h066: out <= 24'hffffff;    10'h0e6: out <= 24'hffffff;    10'h166: out <= 24'h8a6e47;    10'h1e6: out <= 24'h8a6e47;    10'h266: out <= 24'h8a6e47;    10'h2e6: out <= 24'h8a6e47;    10'h366: out <= 24'h8a6e47;    10'h3e6: out <= 24'h000000;
  10'h067: out <= 24'hffffff;    10'h0e7: out <= 24'hffffff;    10'h167: out <= 24'h8a6e47;    10'h1e7: out <= 24'h8a6e47;    10'h267: out <= 24'h404f2c;    10'h2e7: out <= 24'h8a6e47;    10'h367: out <= 24'h404f2c;    10'h3e7: out <= 24'h000000;
  10'h068: out <= 24'hffffff;    10'h0e8: out <= 24'h000000;    10'h168: out <= 24'h8a6e47;    10'h1e8: out <= 24'h8a6e47;    10'h268: out <= 24'h000000;    10'h2e8: out <= 24'h000000;    10'h368: out <= 24'h8a6e47;    10'h3e8: out <= 24'h000000;
  10'h069: out <= 24'hffffff;    10'h0e9: out <= 24'h000000;    10'h169: out <= 24'h8a6e47;    10'h1e9: out <= 24'h000000;    10'h269: out <= 24'hffffff;    10'h2e9: out <= 24'hffffff;    10'h369: out <= 24'h8a6e47;    10'h3e9: out <= 24'h000000;
  10'h06a: out <= 24'hffffff;    10'h0ea: out <= 24'h8a6e47;    10'h16a: out <= 24'h8a6e47;    10'h1ea: out <= 24'hffffff;    10'h26a: out <= 24'hffffff;    10'h2ea: out <= 24'h000000;    10'h36a: out <= 24'h000000;    10'h3ea: out <= 24'h000000;
  10'h06b: out <= 24'hffffff;    10'h0eb: out <= 24'h8a6e47;    10'h16b: out <= 24'h000000;    10'h1eb: out <= 24'hffffff;    10'h26b: out <= 24'hffffff;    10'h2eb: out <= 24'h8a6e47;    10'h36b: out <= 24'hffc18f;    10'h3eb: out <= 24'h000000;
  10'h06c: out <= 24'h000000;    10'h0ec: out <= 24'h8a6e47;    10'h16c: out <= 24'h000000;    10'h1ec: out <= 24'hffffff;    10'h26c: out <= 24'hffffff;    10'h2ec: out <= 24'h8a6e47;    10'h36c: out <= 24'hffc18f;    10'h3ec: out <= 24'h000000;
  10'h06d: out <= 24'h000000;    10'h0ed: out <= 24'h000000;    10'h16d: out <= 24'hffffff;    10'h1ed: out <= 24'hffffff;    10'h26d: out <= 24'h000000;    10'h2ed: out <= 24'h000000;    10'h36d: out <= 24'hffc18f;    10'h3ed: out <= 24'h000000;
  10'h06e: out <= 24'h000000;    10'h0ee: out <= 24'h000000;    10'h16e: out <= 24'hffffff;    10'h1ee: out <= 24'hffffff;    10'h26e: out <= 24'h000000;    10'h2ee: out <= 24'h000000;    10'h36e: out <= 24'hffc18f;    10'h3ee: out <= 24'h000000;
  10'h06f: out <= 24'h000000;    10'h0ef: out <= 24'h000000;    10'h16f: out <= 24'hffffff;    10'h1ef: out <= 24'hffffff;    10'h26f: out <= 24'h000000;    10'h2ef: out <= 24'hffc18f;    10'h36f: out <= 24'hffc18f;    10'h3ef: out <= 24'h000000;
  10'h070: out <= 24'h000000;    10'h0f0: out <= 24'h000000;    10'h170: out <= 24'hffffff;    10'h1f0: out <= 24'hffffff;    10'h270: out <= 24'h000000;    10'h2f0: out <= 24'hffc18f;    10'h370: out <= 24'h886028;    10'h3f0: out <= 24'h000000;
  10'h071: out <= 24'h000000;    10'h0f1: out <= 24'h000000;    10'h171: out <= 24'hffffff;    10'h1f1: out <= 24'hffffff;    10'h271: out <= 24'h000000;    10'h2f1: out <= 24'h000000;    10'h371: out <= 24'h886028;    10'h3f1: out <= 24'h000000;
  10'h072: out <= 24'h000000;    10'h0f2: out <= 24'h000000;    10'h172: out <= 24'hffffff;    10'h1f2: out <= 24'hffffff;    10'h272: out <= 24'h000000;    10'h2f2: out <= 24'h000000;    10'h372: out <= 24'h886028;    10'h3f2: out <= 24'h000000;
  10'h073: out <= 24'h000000;    10'h0f3: out <= 24'h000000;    10'h173: out <= 24'hffffff;    10'h1f3: out <= 24'hffffff;    10'h273: out <= 24'hffffff;    10'h2f3: out <= 24'h404f2c;    10'h373: out <= 24'h886028;    10'h3f3: out <= 24'h000000;
  10'h074: out <= 24'h000000;    10'h0f4: out <= 24'h8a6e47;    10'h174: out <= 24'h000000;    10'h1f4: out <= 24'hffffff;    10'h274: out <= 24'hffffff;    10'h2f4: out <= 24'h8a6e47;    10'h374: out <= 24'hffc18f;    10'h3f4: out <= 24'h000000;
  10'h075: out <= 24'hffffff;    10'h0f5: out <= 24'h8a6e47;    10'h175: out <= 24'h000000;    10'h1f5: out <= 24'hffffff;    10'h275: out <= 24'hffffff;    10'h2f5: out <= 24'h000000;    10'h375: out <= 24'h000000;    10'h3f5: out <= 24'h000000;
  10'h076: out <= 24'hffffff;    10'h0f6: out <= 24'h404f2c;    10'h176: out <= 24'h8a6e47;    10'h1f6: out <= 24'h000000;    10'h276: out <= 24'hffffff;    10'h2f6: out <= 24'hffffff;    10'h376: out <= 24'h8a6e47;    10'h3f6: out <= 24'h000000;
  10'h077: out <= 24'hffffff;    10'h0f7: out <= 24'h000000;    10'h177: out <= 24'h8a6e47;    10'h1f7: out <= 24'h8a6e47;    10'h277: out <= 24'h000000;    10'h2f7: out <= 24'h000000;    10'h377: out <= 24'h404f2c;    10'h3f7: out <= 24'h000000;
  10'h078: out <= 24'hffffff;    10'h0f8: out <= 24'h000000;    10'h178: out <= 24'h8a6e47;    10'h1f8: out <= 24'h8a6e47;    10'h278: out <= 24'h8a6e47;    10'h2f8: out <= 24'h8a6e47;    10'h378: out <= 24'h404f2c;    10'h3f8: out <= 24'h000000;
  10'h079: out <= 24'hffffff;    10'h0f9: out <= 24'hffffff;    10'h179: out <= 24'h8a6e47;    10'h1f9: out <= 24'h8a6e47;    10'h279: out <= 24'h8a6e47;    10'h2f9: out <= 24'h8a6e47;    10'h379: out <= 24'h8a6e47;    10'h3f9: out <= 24'h000000;
  10'h07a: out <= 24'hffffff;    10'h0fa: out <= 24'hffffff;    10'h17a: out <= 24'h8a6e47;    10'h1fa: out <= 24'h8a6e47;    10'h27a: out <= 24'h8a6e47;    10'h2fa: out <= 24'h8a6e47;    10'h37a: out <= 24'h8a6e47;    10'h3fa: out <= 24'h000000;
  10'h07b: out <= 24'hffffff;    10'h0fb: out <= 24'hffffff;    10'h17b: out <= 24'h000000;    10'h1fb: out <= 24'h8a6e47;    10'h27b: out <= 24'h8a6e47;    10'h2fb: out <= 24'h8a6e47;    10'h37b: out <= 24'h404f2c;    10'h3fb: out <= 24'hffffff;
  10'h07c: out <= 24'hffffff;    10'h0fc: out <= 24'hffffff;    10'h17c: out <= 24'hffffff;    10'h1fc: out <= 24'h8a6e47;    10'h27c: out <= 24'h8a6e47;    10'h2fc: out <= 24'h8a6e47;    10'h37c: out <= 24'h404f2c;    10'h3fc: out <= 24'hffffff;
  10'h07d: out <= 24'hffffff;    10'h0fd: out <= 24'hffffff;    10'h17d: out <= 24'hffffff;    10'h1fd: out <= 24'h000000;    10'h27d: out <= 24'h000000;    10'h2fd: out <= 24'h000000;    10'h37d: out <= 24'h000000;    10'h3fd: out <= 24'hffffff;
  10'h07e: out <= 24'hffffff;    10'h0fe: out <= 24'hffffff;    10'h17e: out <= 24'hffffff;    10'h1fe: out <= 24'hffffff;    10'h27e: out <= 24'hffffff;    10'h2fe: out <= 24'hffffff;    10'h37e: out <= 24'hffffff;    10'h3fe: out <= 24'hffffff;
  10'h07f: out <= 24'hffffff;    10'h0ff: out <= 24'hffffff;    10'h17f: out <= 24'hffffff;    10'h1ff: out <= 24'hffffff;    10'h27f: out <= 24'hffffff;    10'h2ff: out <= 24'hffffff;    10'h37f: out <= 24'hffffff;    10'h3ff: out <= 24'hffffff;
	endcase
endmodule
