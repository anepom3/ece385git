// We'll create the MAR module here.
