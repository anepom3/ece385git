// We'll create the IR file here!
