// This file is for the ADDR module!
