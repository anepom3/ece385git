// This is the file for the ADDR2MUX!
